`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/29
// Design Name: 
// Module Name: arbitrate_bpsi
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
// `define FBC_UDP_OFF


module arbitrate_bpsi #(
    parameter                               TCQ                 = 0.1   ,
    parameter        [8*20-1:0]             MFPGA_VERSION       = "PCG1_TimingM_v1.1   "
)(
    // clk & rst
    input    wire                           clk_i                       ,
    input    wire                           rst_i                       ,
    input    wire    [64-1:0]               heartbeat_data_i            ,
    input    wire                           heartbeat_en_i              ,
    input    wire    [64-1:0]               readback_data_i             ,
    input    wire                           readback_vld_i              ,
    input    wire    [64-1:0]               fpga_message_up_data_i      ,
    input    wire                           fpga_message_up_i           ,
    input    wire                           ddr_readback_vld_i          ,
    input    wire                           ddr_readback_last_i         ,
    input    wire    [64-1:0]               ddr_readback_data_i         ,

    // // calibrate voltage. dark current * R
    // input    wire                           FBCi_cali_en_i              ,
    // input    wire    [23:0]                 FBCi_cali_a_i               ,
    // input    wire    [23:0]                 FBCi_cali_b_i               ,
    // input    wire                           FBCr1_cali_en_i             ,
    // input    wire    [23:0]                 FBCr1_cali_a_i              ,
    // input    wire    [23:0]                 FBCr1_cali_b_i              ,
    // input    wire                           FBCr2_cali_en_i             ,
    // input    wire    [23:0]                 FBCr2_cali_a_i              ,
    // input    wire    [23:0]                 FBCr2_cali_b_i              ,
    
    // actual voltage
    input    wire                           FBC_out_fifo_rst_i          ,
    input    wire                           fbc_udp_rate_switch_i       ,
    input    wire                           FBC_out_vld_i               ,
    // input    wire                           FBCi_out_en_i               ,
    input    wire    [23:0]                 FBCi_out_a_i                ,
    input    wire    [23:0]                 FBCi_out_b_i                ,
    // input    wire                           FBCr1_out_en_i              ,
    input    wire    [23:0]                 FBCr1_out_a_i               ,
    input    wire    [23:0]                 FBCr1_out_b_i               ,
    // input    wire                           FBCr2_out_en_i              ,
    input    wire    [23:0]                 FBCr2_out_a_i               ,
    input    wire    [23:0]                 FBCr2_out_b_i               ,
    // Enocde
    input    wire    [32-1:0]               encode_w_i                  ,
    input    wire    [32-1:0]               encode_x_i                  ,

    // background voltage. dark current * R
    input    wire                           FBCi_bg_en_i                ,
    input    wire    [23:0]                 FBCi_bg_a_i                 ,
    input    wire    [23:0]                 FBCi_bg_b_i                 ,
    input    wire                           FBCr1_bg_en_i               ,
    input    wire    [23:0]                 FBCr1_bg_a_i                ,
    input    wire    [23:0]                 FBCr1_bg_b_i                ,
    input    wire                           FBCr2_bg_en_i               ,
    input    wire    [23:0]                 FBCr2_bg_a_i                ,
    input    wire    [23:0]                 FBCr2_bg_b_i                ,

    input    wire                           quad_sensor_data_en_i       ,
    input    wire    [96-1:0]               quad_sensor_data_i          ,
    input    wire                           quad_sensor_bg_data_en_i    ,
    input    wire    [96-1:0]               quad_sensor_bg_data_i       ,

    input    wire                           motor_data_in_en_i          , // Uop en
    input    wire    [15:0]                 motor_data_in_i             , // Uop to motor
    input    wire    [15:0]                 motor_data_out_i            , // Ufeed
    
    input    wire    [8-1:0]                laser_rx_data_i             ,
    input    wire                           laser_rx_vld_i              ,
    input    wire                           laser_rx_last_i             ,

    input    wire                           spi_slave0_ack_rst_i        ,
    input    wire                           spi_slave0_ack_vld_i        ,
    input    wire                           spi_slave0_ack_last_i       ,
    input    wire    [32-1:0]               spi_slave0_ack_data_i       ,
    input    wire                           spi_slave1_ack_rst_i        ,
    input    wire                           spi_slave1_ack_vld_i        ,
    input    wire                           spi_slave1_ack_last_i       ,
    input    wire    [32-1:0]               spi_slave1_ack_data_i       ,
    input    wire                           spi_slave2_ack_rst_i        ,
    input    wire                           spi_slave2_ack_vld_i        ,
    input    wire                           spi_slave2_ack_last_i       ,
    input    wire    [32-1:0]               spi_slave2_ack_data_i       ,

    // read mfpga version
    input    wire                           rd_mfpga_version_i          ,

    // eds error row
    input    wire                           eds_error_vld_i             ,
    input    wire   [16-1:0]                eds_error_data_i            ,
    // slave comm
    input    wire                           slave_tx_ack_i              ,
    output   wire                           slave_tx_byte_num_en_o      ,
    output   wire   [15:0]                  slave_tx_byte_num_o         ,
    output   wire                           slave_tx_byte_en_o          ,
    output   wire   [ 7:0]                  slave_tx_byte_o             

);


//////////////////////////////////////////////////////////////////////////////////
// *********** Define Parameter Signal
//>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
localparam          [16-1:0]                FBC_ACTUAL_TYPE             = 'h010F;
localparam          [11-1:0]                FBC_ACTUAL_DATA_NUM         = 'd30;
localparam          [16-1:0]                FBC_ACTUAL_BYTE_NUM         = FBC_ACTUAL_DATA_NUM * 18 + 2 + FBC_ACTUAL_DATA_NUM*8;

localparam          [16-1:0]                FBC_VOL_TYPE                = 'h010B;
localparam          [11-1:0]                FBC_VOL_DATA_NUM            = 'd10;
localparam          [16-1:0]                FBC_VOL_BYTE_NUM            = FBC_VOL_DATA_NUM * 4 + 2;

localparam          [16-1:0]                FBC_BG_CALI_TYPE            = 'h0115;
localparam          [16-1:0]                FBC_BG_CALI_NUM             = 'd21;

localparam          [16-1:0]                LASER_UART_TYPE             = 'h0122;

localparam          [16-1:0]                SPI_SLAVE_ACK_TYPE          = 'h0123;

localparam          [16-1:0]                MFPGA_VERSION_TYPE          = 'h0100;
localparam          [16-1:0]                MFPGA_VERSION_NUM           = 'd22;

localparam          [16-1:0]                READBACK_TYPE               = 'h0200;
localparam          [16-1:0]                READBACK_NUM                = 'd10;

localparam          [16-1:0]                HEARTBEAT_TYPE              = 'h0350;
localparam          [16-1:0]                HEARTBEAT_NUM               = 'd10;

localparam          [16-1:0]                FPGA_ACT_MESS_TYPE          = 'h0340;
localparam          [16-1:0]                FPGA_ACT_MESS_NUM           = 'd10;

localparam          [16-1:0]                DDR_READBACK_TYPE           = 'h035E;
// localparam          [16-1:0]                DDR_READBACK_NUM            = 'd128;  // 128*64 = 1024*8

localparam          [16-1:0]                QUAD_SENSOR_TYPE            = 'h0332;
localparam          [16-1:0]                QUAD_SENSOR_NUM             = FBC_ACTUAL_DATA_NUM * 12 + 2 + FBC_ACTUAL_DATA_NUM*8;

localparam          [16-1:0]                EDS_ERROR_TYPE              = 'h0360;
localparam                                  ARBITRATE_NUM               = 14;    // control arbitrate channel
genvar i;
//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<

//////////////////////////////////////////////////////////////////////////////////
// *********** Define Register Signal
//>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
// reg                                         FBCi_wr_en_d0               = 'd0;
// reg                                         FBCi_wr_en_d1               = 'd0;
// reg                                         FBCr1_wr_en_d0              = 'd0;
// reg                                         FBCr1_wr_en_d1              = 'd0;
// reg                                         FBCr2_wr_en_d0              = 'd0;
// reg                                         FBCr2_wr_en_d1              = 'd0;

reg                                         FBC_out_vld_d0              = 'd0;
reg                                         FBC_out_vld_d1              = 'd0;

reg                 [24-1:0]                FBCi_data_b                 = 'd0;
reg                 [24-1:0]                FBCr1_data_b                = 'd0;
reg                 [24-1:0]                FBCr2_data_b                = 'd0;

reg                 [24-1:0]                FBCi_din                    = 'd0;
reg                 [24-1:0]                FBCr1_din                   = 'd0;
reg                 [24-1:0]                FBCr2_din                   = 'd0;

// reg                 [ 7-1:0]                FBCi_cnt                    = 'd0;
// reg                 [ 7-1:0]                FBCr1_cnt                   = 'd0;
// reg                 [ 7-1:0]                FBCr2_cnt                   = 'd0;
reg                 [ 7-1:0]                FBC_src_cnt                 = 'd0;
reg                 [ 7-1:0]                quad_cnt                    = 'd0;

reg                                         FBCi_rd_en                  = 'd0;
reg                                         FBCr1_rd_en                 = 'd0;
reg                                         FBCr2_rd_en                 = 'd0;
reg                                         fbc_encode_rd               = 'd0;


reg                                         fbc_i_full                  = 'd0;
reg                                         fbc_r1_full                 = 'd0;
reg                                         fbc_r2_full                 = 'd0;
reg                                         quad_full                   = 'd0;

reg                                         fbc_vol_wr_en_d0            = 'd0;
reg                                         fbc_vol_wr_en_d1            = 'd0;
reg                 [16-1:0]                fbc_vol_feed_d              = 'd0;
reg                 [16-1:0]                fbc_vol_din                 = 'd0;
reg                 [ 7-1:0]                fbc_vol_cnt                 = 'd0;
reg                                         fbc_vol_rd_en               = 'd0;

reg                 [10-1:0]                laser_rx_cnt                = 'd0;
reg                 [10-1:0]                laser_rx_num                = 'd0;
reg                                         laser_rx_rd_en              = 'd0;

reg                 [ARBITRATE_NUM-1:0]     arbitrate                   = 'd1;
reg                 [ARBITRATE_NUM-1:0]     bpsi_type                   = 'd0;
reg                                         arbitr_result_d0            = 'd0;
reg                                         arbitr_result_d1            = 'd0;

reg                 [160-1:0]               slave_tx_data               = 'd0;

reg                 [11-1:0]                slave_tx_cnt                = 'd0;
reg                 [ 8-1:0]                slave_tx_byte               = 'd0;
reg                                         slave_tx_byte_en            = 'd0;

reg                 [24-1:0]                FBCi_bg_data_a_sync         = 'd0;
reg                 [24-1:0]                FBCi_bg_data_b_sync         = 'd0;
// reg                 [24-1:0]                FBCi_cali_data_a_sync       = 'd0;
// reg                 [24-1:0]                FBCi_cali_data_b_sync       = 'd0;
reg                 [24-1:0]                FBCr1_bg_data_a_sync        = 'd0;
reg                 [24-1:0]                FBCr1_bg_data_b_sync        = 'd0;
// reg                 [24-1:0]                FBCr1_cali_data_a_sync      = 'd0;
// reg                 [24-1:0]                FBCr1_cali_data_b_sync      = 'd0;
reg                 [24-1:0]                FBCr2_bg_data_a_sync        = 'd0;
reg                 [24-1:0]                FBCr2_bg_data_b_sync        = 'd0;
reg                                         quad_sensor_bg_data_en_d    = 'd0;
reg                 [96-1:0]                quad_sensor_bg_data_d       = 'd0;
reg                 [8-1:0]                 bg_time_share               = 'd0;
reg                 [144-1:0]               bg_time_share_data          = 'd0;
reg                 [16-1:0]                slave_tx_byte_num           = 'd0;

reg                                         FBCi_bg_ready               = 'd0;
reg                                         FBCr1_bg_ready              = 'd0;
reg                                         FBCr2_bg_ready              = 'd0;
// reg                                         FBCi_cali_ready             = 'd0;
// reg                                         FBCr2_cali_ready            = 'd0;
reg                                         quad_sensor_rd              = 'd0;


// ddr readback channel
reg                                         ddr_readback_rd             = 'd0;
reg                 [16-1:0]                ddr_readback_cnt            = 'd0;
reg                 [16-1:0]                ddr_readback_num            = 'd0;

// eds error channel
reg                                         eds_error_rd                = 'd0;

reg                 [ 6-1:0]                spi_slave_ack_cnt [2:0] ;
reg                 [ 6-1:0]                spi_slave_ack_num [2:0] ;
reg                                         spi_ack_rd_en     [2:0] ;
//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<



//////////////////////////////////////////////////////////////////////////////////
// *********** Define Wire Signal
//>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
wire                [ARBITRATE_NUM-1:0]     bpsi_en             ;
wire                [ARBITRATE_NUM-1:0]     arbitr_result       ;

wire                                        FBCi_arbitr_en      ;
wire                                        FBCr1_arbitr_en     ;
wire                                        FBCr2_arbitr_en     ;
wire                [24-1:0]                FBCi_dout           ;
wire                [24-1:0]                FBCr1_dout          ;
wire                [24-1:0]                FBCr2_dout          ;
wire                                        FBCi_full           ;
wire                                        FBCi_empty          ;
wire                                        FBCr1_full          ;
wire                                        FBCr1_empty         ;
wire                                        FBCr2_full          ;
wire                                        FBCr2_empty         ;
wire                                        fbc_encode_vld      ;
wire                [64-1:0]                fbc_encode_data     ;

wire                                        fbc_arbitr_en       ;
wire                                        quad_arbitr_en      ;

wire                                        FBC_bg_arbitr_en    ;
wire                                        bg_arbitr_en        ;
// wire                                        FBC_cali_arbitr_en  ;

wire                [16-1:0]                fbc_vol_dout        ;
wire                                        fbc_vol_arbitr_en   ;

wire                                        laser_rx_en         ;
wire                [ 8-1:0]                laser_rx_dout       ;

wire                                        quad_sensor_vld     ;
wire                [96+64-1:0]             quad_sensor_data    ;

wire                                        ddr_readback_vld    ;
wire                [64-1:0]                ddr_readback_data   ;

wire                                        eds_error_vld       ;
wire                [16-1:0]                eds_error_data      ;

wire                                        spi_slave_ack_en [3:0];
wire                [32-1:0]                spi_ack_rd_dout  [3:0];
wire                                        spi_ack_full     [3:0];
wire                                        spi_ack_empty    [3:0];

//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<





//////////////////////////////////////////////////////////////////////////////////
// *********** Instance Module
//>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
bpsi_fbc_fifo bpsi_fbci_fifo_inst(
  .clk                      ( clk_i                                 ),
  .srst                     ( rst_i || FBC_out_fifo_rst_i           ),
  .din                      ( FBCi_din                              ),
  .wr_en                    ( FBC_out_vld_d1 || FBC_out_vld_d0      ),
  .rd_en                    ( FBCi_rd_en                            ),
  .dout                     ( FBCi_dout                             ),
  .full                     ( FBCi_full                             ),
  .empty                    ( FBCi_empty                            )
);

bpsi_fbc_fifo bpsi_fbcr1_fifo_inst(
  .clk                      ( clk_i                                 ),
  .srst                     ( rst_i || FBC_out_fifo_rst_i           ),
  .din                      ( FBCr1_din                             ),
  .wr_en                    ( FBC_out_vld_d1 || FBC_out_vld_d0      ),
  .rd_en                    ( FBCr1_rd_en                           ),
  .dout                     ( FBCr1_dout                            ),
  .full                     ( FBCr1_full                            ),
  .empty                    ( FBCr1_empty                           )
);

bpsi_fbc_fifo bpsi_fbcr2_fifo_inst(
  .clk                      ( clk_i                                 ),
  .srst                     ( rst_i || FBC_out_fifo_rst_i           ),
  .din                      ( FBCr2_din                             ),
  .wr_en                    ( FBC_out_vld_d1 || FBC_out_vld_d0      ),
  .rd_en                    ( FBCr2_rd_en                           ),
  .dout                     ( FBCr2_dout                            ),
  .full                     ( FBCr2_full                            ),
  .empty                    ( FBCr2_empty                           )
);

xpm_sync_fifo #(
    .ECC_MODE               ( "no_ecc"                              ),
    .FIFO_MEMORY_TYPE       ( "block"                               ), // "auto" "block" "distributed"
    .READ_MODE              ( "fwft"                                ),
    .FIFO_WRITE_DEPTH       ( 256                                   ),
    .WRITE_DATA_WIDTH       ( 64                                    ),
    .READ_DATA_WIDTH        ( 64                                    ),
    .USE_ADV_FEATURES       ( "1808"                                )
)u_xpm_sync_fifo (
    .wr_clk_i               ( clk_i                                 ),
    .rst_i                  ( rst_i || FBC_out_fifo_rst_i           ), // synchronous to wr_clk
    .wr_en_i                ( FBCr2_out_en_i                        ),
    .wr_data_i              ( {encode_w_i,encode_x_i}               ),

    .rd_en_i                ( fbc_encode_rd                         ),
    .fifo_rd_vld_o          ( fbc_encode_vld                        ),
    .fifo_rd_data_o         ( fbc_encode_data                       )
);

xpm_sync_fifo #(
    .ECC_MODE               ( "no_ecc"                              ),
    .FIFO_MEMORY_TYPE       ( "block"                               ), // "auto" "block" "distributed"
    .READ_MODE              ( "fwft"                                ),
    .FIFO_WRITE_DEPTH       ( 256                                   ),
    .WRITE_DATA_WIDTH       ( 96+64                                 ),
    .READ_DATA_WIDTH        ( 96+64                                 ),
    .USE_ADV_FEATURES       ( "1808"                                )
)quad_sensor_fifo (
    .wr_clk_i               ( clk_i                                 ),
    .rst_i                  ( rst_i || FBC_out_fifo_rst_i           ), // synchronous to wr_clk
    .wr_en_i                ( quad_sensor_data_en_i                 ),
    .wr_data_i              ( {quad_sensor_data_i,encode_w_i,encode_x_i}),

    .rd_en_i                ( quad_sensor_rd                        ),
    .fifo_rd_vld_o          ( quad_sensor_vld                       ),
    .fifo_rd_data_o         ( quad_sensor_data                      )
);

fbc_voltage_fifo fbc_voltage_fifo_inst(
  .clk                      ( clk_i                                 ),
  .srst                     ( rst_i                                 ),
  .din                      ( fbc_vol_din                           ),
  .wr_en                    ( fbc_vol_wr_en_d1 || fbc_vol_wr_en_d0  ),
  .rd_en                    ( fbc_vol_rd_en                         ),
  .dout                     ( fbc_vol_dout                          ),
  .full                     ( fbc_vol_full                          ),
  .empty                    ( fbc_vol_empty                         )
);

laser_rx_fifo laser_rx_fifo_inst(
    .clk                    ( clk_i                                 ),
    .srst                   ( rst_i                                 ),
    .din                    ( laser_rx_data_i                       ),
    .wr_en                  ( laser_rx_vld_i                        ),
    .rd_en                  ( laser_rx_rd_en                        ),
    .dout                   ( laser_rx_dout                         ),
    .full                   ( laser_rx_full                         ),
    .empty                  ( laser_rx_empty                        )
);

generate
    for (i = 0; i<3; i=i+1) begin
        spi_slave_ack_fifo spi_slave_ack_fifo_inst(
            .clk            ( clk_i                                 ),
            .srst           ( rst_i                                 ),
            .din            ( spi_slave_ack_data[i]                 ),
            .wr_en          ( spi_slave_ack_vld[i]                  ),
            .rd_en          ( spi_ack_rd_en[i]                      ),
            .dout           ( spi_ack_rd_dout[i]                    ),
            .full           ( spi_ack_full[i]                       ),
            .empty          ( spi_ack_empty[i]                      )
        );
    end
endgenerate

xpm_sync_fifo #(
    .ECC_MODE               ( "no_ecc"                              ),
    .FIFO_MEMORY_TYPE       ( "block"                               ), // "auto" "block" "distributed"
    .READ_MODE              ( "fwft"                                ),
    .FIFO_WRITE_DEPTH       ( 256                                   ),
    .WRITE_DATA_WIDTH       ( 64                                    ),
    .READ_DATA_WIDTH        ( 64                                    ),
    .USE_ADV_FEATURES       ( "1808"                                )
)ddr_readback_inst (
    .wr_clk_i               ( clk_i                                 ),
    .rst_i                  ( rst_i                                 ), // synchronous to wr_clk
    .wr_en_i                ( ddr_readback_vld_i                    ),
    .wr_data_i              ( ddr_readback_data_i                   ),

    .rd_en_i                ( ddr_readback_rd                       ),
    .fifo_rd_vld_o          ( ddr_readback_vld                      ),
    .fifo_rd_data_o         ( ddr_readback_data                     )
);

xpm_sync_fifo #(
    .ECC_MODE               ( "no_ecc"                              ),
    .FIFO_MEMORY_TYPE       ( "block"                               ), // "auto" "block" "distributed"
    .READ_MODE              ( "fwft"                                ),
    .FIFO_WRITE_DEPTH       ( 2048                                  ),
    .WRITE_DATA_WIDTH       ( 16                                    ),
    .READ_DATA_WIDTH        ( 16                                    ),
    .USE_ADV_FEATURES       ( "1808"                                )
)eds_error_row_inst (
    .wr_clk_i               ( clk_i                                 ),
    .rst_i                  ( rst_i                                 ), // synchronous to wr_clk
    .wr_en_i                ( eds_error_vld_i                       ),
    .wr_data_i              ( eds_error_data_i                      ),

    .rd_en_i                ( eds_error_rd                          ),
    .fifo_rd_vld_o          ( eds_error_vld                         ),
    .fifo_rd_data_o         ( eds_error_data                        )
);

//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<


//////////////////////////////////////////////////////////////////////////////////
// *********** Logic Design
//>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>>
// FBCi,FBCr1,FBCr2 data ready. 
// generate a transmission every 100 times.
// fifo width is 3byte,twice write en,for save resources.
always @(posedge clk_i) FBC_out_vld_d0   <= #TCQ FBC_out_vld_i;
always @(posedge clk_i) FBC_out_vld_d1   <= #TCQ FBC_out_vld_d0;

always @(posedge clk_i) FBCi_data_b     <= #TCQ FBCi_out_b_i;
always @(posedge clk_i) FBCr1_data_b    <= #TCQ FBCr1_out_b_i;
always @(posedge clk_i) FBCr2_data_b    <= #TCQ FBCr2_out_b_i;

always @(posedge clk_i) begin
    if(FBC_out_vld_i)begin
        FBCi_din  <= #TCQ FBCi_out_a_i;
        FBCr1_din <= #TCQ FBCr1_out_a_i;
        FBCr2_din <= #TCQ FBCr2_out_a_i;
    end
    else if(FBC_out_vld_d0)begin
        FBCi_din  <= #TCQ FBCi_data_b;
        FBCr1_din <= #TCQ FBCr1_data_b;
        FBCr2_din <= #TCQ FBCr2_data_b;
    end
end

always @(posedge clk_i) begin
    if(rst_i || FBC_out_fifo_rst_i)
        FBC_src_cnt <= #TCQ 'd0;
    else if(FBC_out_vld_d1)begin
        if(FBC_src_cnt == FBC_ACTUAL_DATA_NUM - 1)
            FBC_src_cnt <= #TCQ 'd0;
        else
            FBC_src_cnt <= #TCQ FBC_src_cnt + 1;
    end
end

assign fbc_arbitr_en = (FBC_src_cnt == FBC_ACTUAL_DATA_NUM - 1) && FBC_out_vld_d1;
// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate fbc_sensor enable end

// qbd quad sensor data ready
always @(posedge clk_i) begin
    if(rst_i || FBC_out_fifo_rst_i)
        quad_cnt <= #TCQ 'd0;
    else if(quad_sensor_data_en_i)begin
        if(quad_cnt == FBC_ACTUAL_DATA_NUM - 1)
            quad_cnt <= #TCQ 'd0;
        else 
            quad_cnt <= #TCQ quad_cnt + 1;
    end
end

assign quad_arbitr_en = (quad_cnt == FBC_ACTUAL_DATA_NUM - 1) && quad_sensor_data_en_i;

// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate quad sensor enable end

// fbc_background_voltage and fbc_cali_position data ready.
always @(posedge clk_i) begin
    if(FBCi_bg_en_i)begin
        FBCi_bg_data_a_sync <= #TCQ FBCi_bg_a_i;
        FBCi_bg_data_b_sync <= #TCQ FBCi_bg_b_i;
    end
end

always @(posedge clk_i) begin
    if(FBCr1_bg_en_i)begin
        FBCr1_bg_data_a_sync <= #TCQ FBCr1_bg_a_i;
        FBCr1_bg_data_b_sync <= #TCQ FBCr1_bg_b_i;
    end 
end

always @(posedge clk_i) begin
    if(FBCr2_bg_en_i)begin
        FBCr2_bg_data_a_sync <= #TCQ FBCr2_bg_a_i;
        FBCr2_bg_data_b_sync <= #TCQ FBCr2_bg_b_i;
    end
end

always @(posedge clk_i) begin
    quad_sensor_bg_data_en_d <= #TCQ quad_sensor_bg_data_en_i;
    if(quad_sensor_bg_data_en_i) quad_sensor_bg_data_d <= #TCQ quad_sensor_bg_data_i;
end

always @(posedge clk_i) begin
    if(FBCi_bg_en_i)            FBCi_bg_ready <= #TCQ 'd1;
    else if(FBC_bg_arbitr_en)   FBCi_bg_ready <= #TCQ 'd0;
    
    if(FBCr1_bg_en_i)           FBCr1_bg_ready <= #TCQ 'd1;
    else if(FBC_bg_arbitr_en)   FBCr1_bg_ready <= #TCQ 'd0;
    
    if(FBCr2_bg_en_i)           FBCr2_bg_ready <= #TCQ 'd1;
    else if(FBC_bg_arbitr_en)   FBCr2_bg_ready <= #TCQ 'd0;
end
assign FBC_bg_arbitr_en = (FBCi_bg_ready && FBCr1_bg_ready && FBCr2_bg_ready);

assign bg_arbitr_en = FBC_bg_arbitr_en ||  quad_sensor_bg_data_en_d;

always @(posedge clk_i) begin
    if(FBC_bg_arbitr_en)
        bg_time_share <= #TCQ 'd2;
    else if(quad_sensor_bg_data_en_d)
        bg_time_share <= #TCQ 'd1;
end
always @(posedge clk_i) begin
    if(FBC_bg_arbitr_en)
        bg_time_share_data <= #TCQ { FBCi_bg_data_a_sync[23:0],FBCi_bg_data_b_sync[23:0]
                                    ,FBCr1_bg_data_a_sync[23:0],FBCr1_bg_data_b_sync[23:0]
                                    ,FBCr2_bg_data_a_sync[23:0],FBCr2_bg_data_b_sync[23:0]};
    else if(quad_sensor_bg_data_en_d)
        bg_time_share_data <= #TCQ {quad_sensor_bg_data_d,48'd0};
end

// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate fbc_background and fbc_calibration enable end

// FBC_Uop FBC_Ufeed data ready. 
// generate a transmission every 10 times.
// fifo width is 2byte,twice write en,for save resources.
always @(posedge clk_i) fbc_vol_wr_en_d0 <= #TCQ motor_data_in_en_i;
always @(posedge clk_i) fbc_vol_wr_en_d1 <= #TCQ fbc_vol_wr_en_d0;

always @(posedge clk_i) fbc_vol_feed_d <= #TCQ motor_data_out_i;
always @(posedge clk_i) begin
    if(motor_data_in_en_i)
        fbc_vol_din <= #TCQ motor_data_in_i;
    else if(fbc_vol_wr_en_d0)
        fbc_vol_din <= #TCQ fbc_vol_feed_d;
end

always @(posedge clk_i) begin
    if(fbc_vol_wr_en_d1)begin
        if(fbc_vol_cnt == FBC_VOL_DATA_NUM - 1)
            fbc_vol_cnt <= #TCQ 'd0;
        else 
            fbc_vol_cnt <= #TCQ fbc_vol_cnt + 1;
    end
end

assign fbc_vol_arbitr_en = (fbc_vol_cnt == FBC_VOL_DATA_NUM - 1) && fbc_vol_wr_en_d1;
// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate fbc_uop and fbc_ufeed enable end 

// generate laser_rx enable
// when laser_rx_last, upload LASER_RX_NUM and sync enable. 
always @(posedge clk_i) begin
    if(laser_rx_vld_i && ~laser_rx_last_i)
        laser_rx_cnt <= #TCQ laser_rx_cnt + 1;
    else if(laser_rx_last_i)
        laser_rx_cnt <= #TCQ 'd0;
end

always @(posedge clk_i) begin
    if(laser_rx_last_i)
        laser_rx_num <= #TCQ laser_rx_cnt + 1;
end

assign laser_rx_en = laser_rx_vld_i && laser_rx_last_i;

// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate laser_rx enable end
wire            spi_slave_ack_vld  [3:0];
wire            spi_slave_ack_last [3:0];
wire [32-1:0]   spi_slave_ack_data [3:0];

assign  spi_slave_ack_vld [0] = spi_slave0_ack_vld_i ;
assign  spi_slave_ack_last[0] = spi_slave0_ack_last_i;
assign  spi_slave_ack_data[0] = spi_slave0_ack_data_i;
assign  spi_slave_ack_vld [1] = spi_slave1_ack_vld_i ;
assign  spi_slave_ack_last[1] = spi_slave1_ack_last_i;
assign  spi_slave_ack_data[1] = spi_slave1_ack_data_i;
assign  spi_slave_ack_vld [2] = spi_slave2_ack_vld_i ;
assign  spi_slave_ack_last[2] = spi_slave2_ack_last_i;
assign  spi_slave_ack_data[2] = spi_slave2_ack_data_i;
// assign  spi_slave_ack_vld [3] = spi_slave3_ack_vld_i ;
// assign  spi_slave_ack_last[3] = spi_slave3_ack_last_i;
// assign  spi_slave_ack_data[3] = spi_slave3_ack_data_i;

// generate new arbitrate enable
// generate spi slave ack enable, from PMT board
generate
    for (i=0;i<3;i=i+1) begin
        always @(posedge clk_i) begin
            if(rst_i)
                spi_slave_ack_cnt[i] <= #TCQ 'd0;
            else if(spi_slave_ack_vld[i] && ~spi_slave_ack_last[i])
                spi_slave_ack_cnt[i] <= #TCQ spi_slave_ack_cnt[i] + 1;
            else if(spi_slave_ack_last[i])
                spi_slave_ack_cnt[i] <= #TCQ 'd0;
        end
        
        always @(posedge clk_i) begin
            if(spi_slave_ack_last[i])
                spi_slave_ack_num[i] <= #TCQ spi_slave_ack_cnt[i] + 1;
        end
        
        assign spi_slave_ack_en[i] = spi_slave_ack_last[i];
    end
endgenerate

// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate new_arbitrate enable end

wire          ddr_readback_irq ;
// generate new arbitrate enable
// ddr readback
// always @(posedge clk_i) begin
//     if(rst_i)
//         ddr_readback_cnt <= #TCQ 'd0;
//     else if(ddr_readback_last_i)
//         ddr_readback_cnt <= #TCQ 'd0;
//     else if(ddr_readback_vld_i)
//         ddr_readback_cnt <= #TCQ ddr_readback_cnt + 1;
// end

// always @(posedge clk_i) begin
//     if(ddr_readback_last_i)
//         ddr_readback_num <= #TCQ ddr_readback_cnt + 1;
// end

assign ddr_readback_irq = ddr_readback_last_i;

// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< generate ddr readback enable end

wire [2-1:0] eds_error_action ;
assign eds_error_action = {eds_error_vld_i,eds_error_rd};

reg [12-1:0] eds_error_cnt = 'd0;
always @(posedge clk_i) begin
    if(eds_error_action==2'b10)
        eds_error_cnt <= #TCQ eds_error_cnt + 1;
    else if(eds_error_action==2'b01)
        eds_error_cnt <= #TCQ eds_error_cnt - 1;
    else
        eds_error_cnt <= #TCQ eds_error_cnt;
end

reg eds_error_irq = 'd0;
always @(posedge clk_i) begin
    eds_error_irq <= #TCQ (~arbitr_result[13]) && (eds_error_cnt >= 511);
end

// generate arbitrate enable , alwaye modify when arbitrate channel add.
assign bpsi_en          = {  
                             eds_error_irq
                            ,ddr_readback_irq
                            ,fpga_message_up_i
                            ,heartbeat_en_i
                            ,readback_vld_i
                            ,rd_mfpga_version_i
                            ,spi_slave_ack_en[2]
                            ,spi_slave_ack_en[1]
                            ,spi_slave_ack_en[0]
                            ,laser_rx_en
                            ,fbc_vol_arbitr_en
                            ,quad_arbitr_en
                            ,bg_arbitr_en
                            ,fbc_arbitr_en };

assign arbitr_result    = bpsi_type & arbitrate;

// arbitr trigger
generate
    for(i=0;i<ARBITRATE_NUM;i=i+1)begin
        always @(posedge clk_i) begin
            if(bpsi_en[i])
                bpsi_type[i] <= #TCQ 1'b1;
            else if(slave_tx_ack_i && arbitr_result[i])
                bpsi_type[i] <= #TCQ 1'b0;
        end
    end
endgenerate

// check arbitr
always @(posedge clk_i) begin
    if(rst_i)
        arbitrate <= #TCQ 'd1;
    else if(arbitr_result=='d0)
        arbitrate <= #TCQ {arbitrate[ARBITRATE_NUM-2:0],arbitrate[ARBITRATE_NUM-1]};
    else 
        arbitrate <= #TCQ arbitrate;
end
// <<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<< arbitrate control , no need to change

// with arbitrate number change
always @(posedge clk_i) begin
    if(arbitr_result[1])
        slave_tx_data <= #TCQ {8'd0,bg_time_share[7:0] ,bg_time_share_data};

    if(arbitr_result[8])
        slave_tx_data <= #TCQ MFPGA_VERSION;
end

// FBC sensor byte control
reg [2:0] fbc_cnt  = 'd5;
reg [1:0] fbc_byte_cnt = 'd2;
reg [11-1:0] fbc_tx_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[0] && fbc_tx_cnt>='d1 && (fbc_tx_cnt<FBC_ACTUAL_DATA_NUM + 2))begin
        if(fbc_byte_cnt=='d2 && fbc_cnt=='d5)begin
            fbc_byte_cnt <= #TCQ 'd0;
            fbc_cnt      <= #TCQ 'd0;
        end
        else if(fbc_byte_cnt=='d2)begin
            fbc_byte_cnt <= #TCQ 'd0;
            fbc_cnt      <= #TCQ fbc_cnt + 1;
        end
        else begin
            fbc_byte_cnt <= #TCQ fbc_byte_cnt + 1;
            fbc_cnt      <= #TCQ fbc_cnt;
        end
    end
    else begin
        fbc_byte_cnt <= #TCQ 'd2;
        fbc_cnt      <= #TCQ 'd5;
    end
end

reg [2:0] fbc_encode_byte_cnt  = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[0] && (fbc_tx_cnt>=FBC_ACTUAL_DATA_NUM + 2))begin
        if(fbc_encode_byte_cnt=='d7)
            fbc_encode_byte_cnt <= #TCQ 'd0;
        else 
            fbc_encode_byte_cnt <= #TCQ fbc_encode_byte_cnt + 1;
    end
    else 
        fbc_encode_byte_cnt <= #TCQ 'd0;
end

always @(posedge clk_i) begin
    if(arbitr_result[0])begin
        if(fbc_tx_cnt<FBC_ACTUAL_DATA_NUM + 2 && fbc_cnt=='d5 && fbc_byte_cnt=='d2)begin
            fbc_tx_cnt <= #TCQ fbc_tx_cnt + 1;
        end
        else if(fbc_tx_cnt>=FBC_ACTUAL_DATA_NUM + 2 && fbc_encode_byte_cnt=='d7)begin
            fbc_tx_cnt <= #TCQ fbc_tx_cnt + 1;
        end
    end
    else begin
        fbc_tx_cnt <= #TCQ 'd0;
    end
end

// spi ack
reg [2-1:0] spi_byte_cnt = 'd0;
reg [6-1:0] spi_ack_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[5])begin
        if(spi_ack_cnt < 'd2)begin
            spi_ack_cnt  <= #TCQ spi_ack_cnt + 1;
            spi_byte_cnt <= #TCQ 'd0;
        end
        else if(spi_ack_cnt < spi_slave_ack_num[0]+2) begin
            spi_ack_cnt  <= #TCQ (spi_byte_cnt=='d3) ? spi_ack_cnt + 1 : spi_ack_cnt;
            spi_byte_cnt <= #TCQ (spi_byte_cnt=='d3) ? 'd0 : spi_byte_cnt + 1;
        end
        else begin
            spi_ack_cnt  <= #TCQ spi_slave_ack_num[0]+3;
            spi_byte_cnt <= #TCQ 'd0;
        end
    end
    else if(arbitr_result[6])begin
        if(spi_ack_cnt < 'd2)begin
            spi_ack_cnt  <= #TCQ spi_ack_cnt + 1;
            spi_byte_cnt <= #TCQ 'd0;
        end
        else if(spi_ack_cnt < spi_slave_ack_num[1]+2) begin
            spi_ack_cnt  <= #TCQ (spi_byte_cnt=='d3) ? spi_ack_cnt + 1 : spi_ack_cnt;
            spi_byte_cnt <= #TCQ (spi_byte_cnt=='d3) ? 'd0 : spi_byte_cnt + 1;
        end
        else begin
            spi_ack_cnt  <= #TCQ spi_slave_ack_num[1]+3;
            spi_byte_cnt <= #TCQ 'd0;
        end
    end
    else if(arbitr_result[7])begin
        if(spi_ack_cnt < 'd2)begin
            spi_ack_cnt  <= #TCQ spi_ack_cnt + 1;
            spi_byte_cnt <= #TCQ 'd0;
        end
        else if(spi_ack_cnt < spi_slave_ack_num[2]+2) begin
            spi_ack_cnt  <= #TCQ (spi_byte_cnt=='d3) ? spi_ack_cnt + 1 : spi_ack_cnt;
            spi_byte_cnt <= #TCQ (spi_byte_cnt=='d3) ? 'd0 : spi_byte_cnt + 1;
        end
        else begin
            spi_ack_cnt  <= #TCQ spi_slave_ack_num[2]+3;
            spi_byte_cnt <= #TCQ 'd0;
        end
    end
    else begin
        spi_ack_cnt <= #TCQ 'd0;
        spi_byte_cnt <= #TCQ 'd0;
    end
end


reg [1:0] byte_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[3])begin
        if(slave_tx_cnt >= 'd2)begin
            byte_cnt <= #TCQ (byte_cnt=='d1) ? 'd0 : (byte_cnt + 1);
        end
    end
    else begin
        byte_cnt <= #TCQ 'd0;
    end
end

always @(posedge clk_i) begin
    if(arbitr_result[1])begin
        if(slave_tx_cnt < FBC_BG_CALI_NUM + 1)
            slave_tx_cnt <= #TCQ slave_tx_cnt + 1;
    end
    else if(arbitr_result[8])begin
        if(slave_tx_cnt < MFPGA_VERSION_NUM + 1)
            slave_tx_cnt <= #TCQ slave_tx_cnt + 1;
    end
    else if(arbitr_result[3])begin
        if(slave_tx_cnt < 'd3)begin
            slave_tx_cnt <= #TCQ slave_tx_cnt + 1;
        end
        else if(slave_tx_cnt < FBC_VOL_DATA_NUM*2+3)begin
            slave_tx_cnt <= #TCQ (byte_cnt=='d0) ? (slave_tx_cnt + 1) : slave_tx_cnt;
        end
    end
    else if(arbitr_result[4])begin
        if(slave_tx_cnt<laser_rx_num+3)
            slave_tx_cnt <= #TCQ slave_tx_cnt + 1;
    end
    else begin
        slave_tx_cnt <= #TCQ 'd0;
    end
end

always @(posedge clk_i) begin
    if((arbitr_result[0]) && (fbc_tx_cnt<FBC_ACTUAL_DATA_NUM + 2) && slave_tx_byte_en && fbc_byte_cnt=='d1)begin
        FBCi_rd_en  <= #TCQ fbc_cnt[2:1]=='b00;
        FBCr1_rd_en <= #TCQ fbc_cnt[2:1]=='b01;
        FBCr2_rd_en <= #TCQ fbc_cnt[2:1]=='b10;
    end
    else begin
        FBCi_rd_en  <= #TCQ 'd0;
        FBCr1_rd_en <= #TCQ 'd0;
        FBCr2_rd_en <= #TCQ 'd0;
    end
end

always @(posedge clk_i) begin
    if((arbitr_result[0]) && (fbc_tx_cnt>=FBC_ACTUAL_DATA_NUM + 2) && slave_tx_byte_en && fbc_encode_byte_cnt=='d6)
        fbc_encode_rd <= #TCQ 'd1;
    else 
        fbc_encode_rd <= #TCQ 'd0;
end

always @(posedge clk_i) begin  // rd_en to slave_tx_byte need 1clk
    if(byte_cnt=='d0 && slave_tx_cnt >= 'd2 && slave_tx_cnt < FBC_VOL_DATA_NUM*2+3)
        fbc_vol_rd_en <= #TCQ (arbitr_result[3]) && slave_tx_byte_en;
    else 
        fbc_vol_rd_en <= #TCQ 'd0;
end

always @(posedge clk_i) begin  // rd_en to slave_tx_byte need 1clk
    if(slave_tx_cnt > 'd0 && slave_tx_cnt < laser_rx_num + 1)
        laser_rx_rd_en <= #TCQ (arbitr_result[4]) && slave_tx_byte_en;
    else 
        laser_rx_rd_en <= #TCQ 'd0;
end

always @(posedge clk_i) begin  // rd_en to slave_tx_byte need 1clk
    if(spi_ack_cnt > 'd1 && spi_byte_cnt =='d2)begin
        spi_ack_rd_en[0] <= #TCQ (arbitr_result[5]) && slave_tx_byte_en;
        spi_ack_rd_en[1] <= #TCQ (arbitr_result[6]) && slave_tx_byte_en;
        spi_ack_rd_en[2] <= #TCQ (arbitr_result[7]) && slave_tx_byte_en;
    end
    else begin
        spi_ack_rd_en[0] <= #TCQ 'd0;
        spi_ack_rd_en[1] <= #TCQ 'd0;
        spi_ack_rd_en[2] <= #TCQ 'd0;
    end
end

reg [3:0] readback_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[9])begin
        if(readback_cnt < READBACK_NUM + 1)
            readback_cnt <= #TCQ readback_cnt + 1;
    end
    else 
        readback_cnt <= #TCQ 'd0;
end

reg [3:0] heartbeat_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[10])begin
        if(heartbeat_cnt < HEARTBEAT_NUM + 1)
            heartbeat_cnt <= #TCQ heartbeat_cnt + 1;
    end
    else 
        heartbeat_cnt <= #TCQ 'd0;
end

reg [3:0] fpga_act_mess_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[11])begin
        if(fpga_act_mess_cnt < FPGA_ACT_MESS_NUM + 1)
            fpga_act_mess_cnt <= #TCQ fpga_act_mess_cnt + 1;
    end
    else 
        fpga_act_mess_cnt <= #TCQ 'd0;
end

reg [3-1:0] ddr_readback_tx_byte_cnt = 'd7;
reg [16-1:0] ddr_readback_tx_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[12] && (ddr_readback_tx_cnt >= 'd1) && (ddr_readback_tx_cnt < 'd128 + 2))begin
        if(ddr_readback_tx_byte_cnt == 'd7)
            ddr_readback_tx_byte_cnt <= #TCQ 'd0;
        else 
            ddr_readback_tx_byte_cnt <= #TCQ ddr_readback_tx_byte_cnt + 1;
    end
    else 
        ddr_readback_tx_byte_cnt <= #TCQ 'd7;
end

always @(posedge clk_i) begin
    if(arbitr_result[12])begin
        if(ddr_readback_tx_byte_cnt == 'd7)
            ddr_readback_tx_cnt <= #TCQ ddr_readback_tx_cnt + 1;
    end
    else 
        ddr_readback_tx_cnt <= #TCQ 'd0;
end

always @(posedge clk_i) begin
    if((arbitr_result[12]) && (ddr_readback_tx_cnt < 'd128 + 2) && slave_tx_byte_en && (ddr_readback_tx_byte_cnt == 'd6))
        ddr_readback_rd  <= #TCQ 'd1;
    else 
        ddr_readback_rd  <= #TCQ 'd0;
end

reg [2-1:0] eds_error_tx_byte_cnt = 'd1;
reg [16-1:0] eds_error_tx_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[13] && (eds_error_tx_cnt >= 'd1) && (eds_error_tx_cnt < 'd512 + 2))begin
        if(eds_error_tx_byte_cnt == 'd1)
            eds_error_tx_byte_cnt <= #TCQ 'd0;
        else 
            eds_error_tx_byte_cnt <= #TCQ eds_error_tx_byte_cnt + 1;
    end
    else 
        eds_error_tx_byte_cnt <= #TCQ 'd1;
end

always @(posedge clk_i) begin
    if(arbitr_result[13])begin
        if(eds_error_tx_byte_cnt == 'd1)
            eds_error_tx_cnt <= #TCQ eds_error_tx_cnt + 1;
    end
    else 
        eds_error_tx_cnt <= #TCQ 'd0;
end

always @(posedge clk_i) begin
    if((arbitr_result[13]) && (eds_error_tx_cnt < 'd512 + 2) && slave_tx_byte_en && (eds_error_tx_byte_cnt == 'd0))
        eds_error_rd  <= #TCQ 'd1;
    else 
        eds_error_rd  <= #TCQ 'd0;
end


reg [5-1:0] quad_sensor_byte_cnt = 'd19;
reg [16-1:0] quad_sensor_cnt = 'd0;
always @(posedge clk_i) begin
    if(arbitr_result[2] && (quad_sensor_cnt >= 'd1) && (quad_sensor_cnt < FBC_ACTUAL_DATA_NUM + 2))begin
        if(quad_sensor_byte_cnt == 'd19)
            quad_sensor_byte_cnt <= #TCQ 'd0;
        else 
            quad_sensor_byte_cnt <= #TCQ quad_sensor_byte_cnt + 1;
    end
    else 
        quad_sensor_byte_cnt <= #TCQ 'd19;
end

always @(posedge clk_i) begin
    if(arbitr_result[2])begin
        if(quad_sensor_byte_cnt == 'd19)
            quad_sensor_cnt <= #TCQ quad_sensor_cnt + 1;
    end
    else 
        quad_sensor_cnt <= #TCQ 'd0;
end

always @(posedge clk_i) begin
    if((arbitr_result[2]) && (quad_sensor_cnt<FBC_ACTUAL_DATA_NUM + 2) && slave_tx_byte_en && quad_sensor_byte_cnt=='d18)
        quad_sensor_rd  <= #TCQ 'd1;
    else 
        quad_sensor_rd  <= #TCQ 'd0;
end

always @(posedge clk_i) begin
    if(arbitr_result[0])begin
        if(fbc_tx_cnt=='d0)
            slave_tx_byte <= #TCQ FBC_ACTUAL_TYPE[15:8];
        else if(fbc_tx_cnt=='d1)
            slave_tx_byte <= #TCQ FBC_ACTUAL_TYPE[7:0];
        else if(fbc_tx_cnt < FBC_ACTUAL_DATA_NUM + 2)begin
            case(fbc_cnt[2:1])
            'b00 : slave_tx_byte <= #TCQ FBCi_dout[(2-fbc_byte_cnt)*8 +: 8];
            'b01 : slave_tx_byte <= #TCQ FBCr1_dout[(2-fbc_byte_cnt)*8 +: 8];
            'b10 : slave_tx_byte <= #TCQ FBCr2_dout[(2-fbc_byte_cnt)*8 +: 8];
            default : /*default*/;
            endcase
        end
        else begin
            slave_tx_byte <= #TCQ fbc_encode_data[(7-fbc_encode_byte_cnt)*8 +: 8];
        end
    end
    else if((arbitr_result[1]) && slave_tx_cnt < FBC_BG_CALI_NUM)begin
        case(slave_tx_cnt)
            'd0 : slave_tx_byte <= #TCQ FBC_BG_CALI_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ FBC_BG_CALI_TYPE[7:0];
            default: slave_tx_byte <= #TCQ slave_tx_data[(FBC_BG_CALI_NUM - slave_tx_cnt - 1)*8 +: 8];
        endcase
    end
    else if(arbitr_result[2])begin
        case(quad_sensor_cnt)
            'd0 : slave_tx_byte <= #TCQ QUAD_SENSOR_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ QUAD_SENSOR_TYPE[7:0];
            default:slave_tx_byte <= #TCQ quad_sensor_data[(5'd19-quad_sensor_byte_cnt)*8 +: 8];
        endcase
    end
    else if((arbitr_result[8]) && slave_tx_cnt < MFPGA_VERSION_NUM)begin
        case(slave_tx_cnt)
            'd0 : slave_tx_byte <= #TCQ MFPGA_VERSION_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ MFPGA_VERSION_TYPE[7:0];
            default: slave_tx_byte <= #TCQ slave_tx_data[(MFPGA_VERSION_NUM - slave_tx_cnt - 1)*8 +: 8];
        endcase
    end
    else if(arbitr_result[3])begin
        case(slave_tx_cnt)
            'd0 : slave_tx_byte <= #TCQ FBC_VOL_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ FBC_VOL_TYPE[7:0];
            default:slave_tx_byte <= #TCQ fbc_vol_dout[(1-byte_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[4])begin
        case(slave_tx_cnt)
            'd0 : slave_tx_byte <= #TCQ LASER_UART_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ LASER_UART_TYPE[7:0];
            default:slave_tx_byte <= #TCQ laser_rx_dout[0 +: 8];
        endcase
    end
    else if(arbitr_result[5])begin
        case(spi_ack_cnt)
            'd0 : slave_tx_byte <= #TCQ SPI_SLAVE_ACK_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ SPI_SLAVE_ACK_TYPE[7:0];
            default:slave_tx_byte <= #TCQ spi_ack_rd_dout[0][(3-spi_byte_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[6])begin
        case(spi_ack_cnt)
            'd0 : slave_tx_byte <= #TCQ SPI_SLAVE_ACK_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ SPI_SLAVE_ACK_TYPE[7:0];
            default:slave_tx_byte <= #TCQ spi_ack_rd_dout[1][(3-spi_byte_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[7])begin
        case(spi_ack_cnt)
            'd0 : slave_tx_byte <= #TCQ SPI_SLAVE_ACK_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ SPI_SLAVE_ACK_TYPE[7:0];
            default:slave_tx_byte <= #TCQ spi_ack_rd_dout[2][(3-spi_byte_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[9] && readback_cnt<READBACK_NUM)begin
        case(readback_cnt)
            'd0 : slave_tx_byte <= #TCQ READBACK_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ READBACK_TYPE[7:0];
            default:slave_tx_byte <= #TCQ readback_data_i[(4'd9-readback_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[10] && heartbeat_cnt<HEARTBEAT_NUM)begin
        case(heartbeat_cnt)
            'd0 : slave_tx_byte <= #TCQ HEARTBEAT_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ HEARTBEAT_TYPE[7:0];
            default:slave_tx_byte <= #TCQ heartbeat_data_i[(4'd9-heartbeat_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[11] && fpga_act_mess_cnt<FPGA_ACT_MESS_NUM)begin
        case(fpga_act_mess_cnt)
            'd0 : slave_tx_byte <= #TCQ FPGA_ACT_MESS_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ FPGA_ACT_MESS_TYPE[7:0];
            default:slave_tx_byte <= #TCQ fpga_message_up_data_i[(4'd9-fpga_act_mess_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[12])begin
        case(ddr_readback_tx_cnt)
            'd0 : slave_tx_byte <= #TCQ DDR_READBACK_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ DDR_READBACK_TYPE[7:0];
            default:slave_tx_byte <= #TCQ ddr_readback_data[('d7-ddr_readback_tx_byte_cnt)*8 +: 8];
        endcase
    end
    else if(arbitr_result[13])begin
        case(eds_error_tx_cnt)
            'd0 : slave_tx_byte <= #TCQ EDS_ERROR_TYPE[15:8];
            'd1 : slave_tx_byte <= #TCQ EDS_ERROR_TYPE[7:0];
            default:slave_tx_byte <= #TCQ eds_error_data[('d1-eds_error_tx_byte_cnt)*8 +: 8];
        endcase
    end
end

wire fbc_tx_byte_en ;
assign fbc_tx_byte_en = (fbc_tx_cnt>'d0) && (fbc_tx_cnt < FBC_ACTUAL_DATA_NUM + 2 + FBC_ACTUAL_DATA_NUM);
reg fbc_tx_byte_en_d = 'd0;
always @(posedge clk_i) fbc_tx_byte_en_d <= #TCQ fbc_tx_byte_en;

wire quad_tx_byte_en ;
assign quad_tx_byte_en = (quad_sensor_cnt>'d0) && (quad_sensor_cnt < FBC_ACTUAL_DATA_NUM + 2);
reg quad_tx_byte_en_d = 'd0;
always @(posedge clk_i) quad_tx_byte_en_d <= #TCQ quad_tx_byte_en;

wire ddr_readback_tx_byte_en ;
assign ddr_readback_tx_byte_en = (ddr_readback_tx_cnt>'d0) && (ddr_readback_tx_cnt < 'd128 + 2);
reg ddr_readback_tx_byte_en_d = 'd0;
always @(posedge clk_i) ddr_readback_tx_byte_en_d <= #TCQ ddr_readback_tx_byte_en;

wire eds_error_tx_byte_en ;
assign eds_error_tx_byte_en = (eds_error_tx_cnt>'d0) && (eds_error_tx_cnt < 'd512 + 2);
reg eds_error_tx_byte_en_d = 'd0;
always @(posedge clk_i) eds_error_tx_byte_en_d <= #TCQ eds_error_tx_byte_en;

always @(*) begin
    if(arbitr_result[0])
        slave_tx_byte_en = fbc_tx_byte_en_d || fbc_tx_byte_en;
    else if(arbitr_result[1])
        slave_tx_byte_en = (slave_tx_cnt>'d0) && (slave_tx_cnt < FBC_BG_CALI_NUM + 1);
    else if(arbitr_result[2])
        slave_tx_byte_en = quad_tx_byte_en_d || quad_tx_byte_en;
    else if(arbitr_result[8])
        slave_tx_byte_en = (slave_tx_cnt>'d0) && (slave_tx_cnt < MFPGA_VERSION_NUM + 1);
    else if(arbitr_result[3])
        slave_tx_byte_en = (slave_tx_cnt>'d0) && (slave_tx_cnt < FBC_VOL_DATA_NUM*2+3);
    else if(arbitr_result[4])
        slave_tx_byte_en = (slave_tx_cnt>'d0) && (slave_tx_cnt < laser_rx_num + 3);
    else if(arbitr_result[5])
        slave_tx_byte_en = (spi_ack_cnt>'d0) && (spi_ack_cnt < spi_slave_ack_num[0] + 3);
    else if(arbitr_result[6])
        slave_tx_byte_en = (spi_ack_cnt>'d0) && (spi_ack_cnt < spi_slave_ack_num[1] + 3);
    else if(arbitr_result[7])
        slave_tx_byte_en = (spi_ack_cnt>'d0) && (spi_ack_cnt < spi_slave_ack_num[2] + 3);
    else if(arbitr_result[9])
        slave_tx_byte_en = (readback_cnt>'d0) && (readback_cnt < READBACK_NUM + 1);
    else if(arbitr_result[10])
        slave_tx_byte_en = (heartbeat_cnt>'d0) && (heartbeat_cnt < HEARTBEAT_NUM + 1);
    else if(arbitr_result[11])
        slave_tx_byte_en = (fpga_act_mess_cnt>'d0) && (fpga_act_mess_cnt < FPGA_ACT_MESS_NUM + 1);
    else if(arbitr_result[12])
        slave_tx_byte_en = ddr_readback_tx_byte_en_d || ddr_readback_tx_byte_en;
    else if(arbitr_result[13])
        slave_tx_byte_en = eds_error_tx_byte_en_d || eds_error_tx_byte_en;
    else 
        slave_tx_byte_en = 'd0;
end

always @(posedge clk_i) begin
    if(arbitr_result[0])
        slave_tx_byte_num <= #TCQ FBC_ACTUAL_BYTE_NUM;
    if(arbitr_result[1])
        slave_tx_byte_num <= #TCQ FBC_BG_CALI_NUM;
    if(arbitr_result[2])
        slave_tx_byte_num <= #TCQ QUAD_SENSOR_NUM;
    if(arbitr_result[8])
        slave_tx_byte_num <= #TCQ MFPGA_VERSION_NUM;
    if(arbitr_result[3])
        slave_tx_byte_num <= #TCQ FBC_VOL_BYTE_NUM;
    if(arbitr_result[4])
        slave_tx_byte_num <= #TCQ laser_rx_num + 2;
    if(arbitr_result[5])
        slave_tx_byte_num <= #TCQ {spi_slave_ack_num[0][5:0],2'b00} + 'd2;
    if(arbitr_result[6])
        slave_tx_byte_num <= #TCQ {spi_slave_ack_num[1][5:0],2'b00} + 'd2;
    if(arbitr_result[7])
        slave_tx_byte_num <= #TCQ {spi_slave_ack_num[2][5:0],2'b00} + 'd2;
    if(arbitr_result[9])
        slave_tx_byte_num <= #TCQ READBACK_NUM;
    if(arbitr_result[10])
        slave_tx_byte_num <= #TCQ HEARTBEAT_NUM;
    if(arbitr_result[11])
        slave_tx_byte_num <= #TCQ FPGA_ACT_MESS_NUM;
    if(arbitr_result[12])
        slave_tx_byte_num <= #TCQ 'd1026;  // {ddr_readback_num,3'b0} + 2;  // 1026
    if(arbitr_result[13])
        slave_tx_byte_num <= #TCQ 'd1026;
end

always @(posedge clk_i) begin
    arbitr_result_d0 <= #TCQ |arbitr_result;
    arbitr_result_d1 <= #TCQ arbitr_result_d0;
end

assign slave_tx_byte_num_en_o = arbitr_result_d0 && (~arbitr_result_d1);
assign slave_tx_byte_num_o    = slave_tx_byte_num;
assign slave_tx_byte_en_o     = slave_tx_byte_en;
assign slave_tx_byte_o        = slave_tx_byte;
//<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<<


endmodule
